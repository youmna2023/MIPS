module instr_mem          // a synthesisable rom implementation  
 (  
      input     [31:0]     pc,  
      output wire    [31:0]          instruction  
 );  
      wire [4: 0] rom_addr = pc[5: 1];   
      reg [31:0] rom[21:0];  
      initial  
      begin  
                rom[0] <= 32'b00100000000010000000000000100000; //addi $t0, $zero, 32 
                rom[1] <= 32'b00100000000010010000000000110111; //addi $t1, $zero, 55  
                rom[2] <= 32'b00000001000010011000000000100100; //and $s0, $t0, $t1 
                rom[3] <= 32'b00000001000010011000000000100101; //or $s0, $t0, $t1  
                rom[4] <= 32'b10101100000100000000000000000100; //sw $s0, 4($zero)  
                rom[5] <= 32'b00000001000010011001000000100010; //sub $s2, $t0, $t1 
                rom[6] <= 32'b10101100000010000000000000001000; //sw $t0, 8($zero)  
                rom[7] <= 32'b00000001000010011001000000100010; //sub $s2, $t0, $t1   
                rom[8] <= 32'b00010010001100100000000000001001; //beq $s1, $s2, error0  
                rom[9] <= 32'b10001100000100010000000000000100; //lw $s1, 4($zero)  
                rom[10] <= 32'b00110010001100100000000001001000; //andi $s2, $s1, 48   
                rom[11] <= 32'b00010010001100100000000000001001; //beq $s1, $s2, error1  
                rom[12] <= 32'b00000010010100011010000000101010; //slt $s4, $s2, $s1 (Last)  
                rom[13] <= 32'b00000010001000001001000000100000; //add $s2, $s1, $0  
                rom[14] <= 32'b00001100000000000000000000001110; //jal last;  
                rom[15] <= 32'b00100000000010000000000000000000; //addi $t0, $0, 0(error0)
                rom[16] <= 32'b00100000000010010000000000000000; //addi $t1, $0, 0 
                rom[17] <= 32'b00100000000010000000000000000001; //addi $t0, $0, 1(error1);
                rom[18] <= 32'b00100000000010010000000000000001; //addi $t1, $0, 1 ;
                rom[19] <= 32'b00110100000010000000000000000000; //ori $t0, $0, 0(error0)
                rom[20] <= 32'b00001000000000000000000000011111; //j EXIT;
      end 
      assign instruction = (pc[31:0] != 0 )? pc[31:0]:32'b0;
 endmodule
